/*
 * Module Name: mod_sub
 * Author(s): Jessica Buentipo
 * Target: FIPS 203 (ML-KEM / Kyber)
 *
 * Description:
 */

module mod_sub(

);

endmodule
