/*
 * Module Name: poly_mul_ntt
 * Author: Kiet Le
 * Description:
 */

module poly_mul_ntt (

);

endmodule
